`include "common.vh"

module MyDesign(
// System signals
  input wire reset_n,
  input wire clk,

// Control signals
  input wire dut_valid,
  output wire dut_ready,

// Input SRAM interface
  output wire dut__tb__sram_input_write_enable,
  output wire [`SRAM_ADDR_RANGE] dut__tb__sram_input_write_address,
  output wire [`SRAM_DATA_RANGE] dut__tb__sram_input_write_data,
  output wire [`SRAM_ADDR_RANGE] dut__tb__sram_input_read_address,
  input  wire [`SRAM_DATA_RANGE] tb__dut__sram_input_read_data,

// Weight SRAM interface
  output wire dut__tb__sram_weight_write_enable,
  output wire [`SRAM_ADDR_RANGE] dut__tb__sram_weight_write_address,
  output wire [`SRAM_DATA_RANGE] dut__tb__sram_weight_write_data,
  output wire [`SRAM_ADDR_RANGE] dut__tb__sram_weight_read_address,
  input  wire [`SRAM_DATA_RANGE] tb__dut__sram_weight_read_data,

// Result SRAM interface
  output wire dut__tb__sram_result_write_enable,
  output wire [`SRAM_ADDR_RANGE] dut__tb__sram_result_write_address,
  output wire [`SRAM_DATA_RANGE] dut__tb__sram_result_write_data,
  output wire [`SRAM_ADDR_RANGE] dut__tb__sram_result_read_address,
  input  wire [`SRAM_DATA_RANGE] tb__dut__sram_result_read_data
);


reg [`SRAM_DATA_RANGE] previous_value;     // register to store accumulated value
wire[`SRAM_DATA_RANGE] current_result;
wire[`SRAM_DATA_RANGE] mac_result_z;
reg[`SRAM_DATA_RANGE] computed_result_reg;
wire[`SRAM_DATA_RANGE] computed_result_wire;
reg[`SRAM_DATA_RANGE] accumulated_reg;

reg [`SRAM_DATA_RANGE/2] matrixAColumns;       // register to number of memory locations to be read from Sram A and B
reg [`SRAM_DATA_RANGE/2] matrixARows;          // register to number of memory locations to be read from Sram A and B

reg [`SRAM_DATA_RANGE/2 ] matrixBColumns;       // register to number of memory locations to be read from Sram A and B
reg [`SRAM_DATA_RANGE/2] matrixBRows;          // register to number of memory locations to be read from Sram A and B


// Declare intermediate registers  to store the address of values to be read from SRAM A and B.
reg [`SRAM_ADDR_RANGE] dut__tb__sram_input_read_address_reg;
reg [`SRAM_ADDR_RANGE] dut__tb__sram_weight_read_address_reg;
reg [`SRAM_ADDR_RANGE] dut__tb__sram_result_write_address_reg;
reg [`SRAM_DATA_RANGE]dut__tb__sram_result_write_data_reg;
reg [`SRAM_DATA_RANGE] sram_result_write_address_reg;


  reg                           set_dut_ready             ;
  reg                           get_array_size            ;
  reg [1:0]                     read_addr_sel             ;
  reg                           all_element_read_completed;
  reg                           compute_accumulation      ;
  reg                           save_array_size           ;
  reg                           write_enable_sel          ;

  wire  [31:0] sum_w;   // Result from FP_add
  reg   [31:0] sum_r;   // Input A of the FP_add 

reg dut_ready_reg; // register to store current DUT state
reg write_enable;
reg read_enable;
reg compute_complete;
reg read_complete;

reg dut__tb__sram_result_write_enable_reg;
reg dut__tb__sram_weight_write_enable_reg;
reg dut__tb__sram_input_write_enable_reg;

reg [2:0] inst_rnd;



reg [ `SRAM_DATA_RANGE/2 ] matrix_A_read_counter;
reg [ `SRAM_DATA_RANGE/2 ] matrix_A_read_counter_1;
reg [ `SRAM_DATA_RANGE/2 ] matrix_A_read_cycle_counter; // Brows
reg [ `SRAM_DATA_RANGE/2 ] matrix_B_read_cycle_counter; // Arows
reg [ `SRAM_DATA_RANGE/2 ] matrix_B_read_counter_1;
reg [ `SRAM_DATA_RANGE/2 ] matrix_B_read_counter_2;
reg [`SRAM_DATA_RANGE] global_read_cycle_counter;
reg [`SRAM_DATA_RANGE] matrixBReadLimit;
reg [`SRAM_DATA_RANGE] numOfReads;
reg [`SRAM_DATA_RANGE ] matrix_C_result_write_address_reg;
reg [`SRAM_DATA_RANGE ]    matrix_A_address;
 reg [`SRAM_DATA_RANGE ]   matrix_A_row_counter;
 reg [`SRAM_DATA_RANGE ]   matrix_A_col_counter;
 reg [`SRAM_DATA_RANGE ]   matrix_B_row_repeat_counter;



 typedef enum bit[2:0] {
    IDLE                              = 3'd0, 
    READ_SRAM_ZERO_ADDR               = 3'd1,   
    READ_SRAM_FIRST_ARRAY_ELEMENT     = 3'd2,   
    READ_SRAM_2_N_ARRAY              = 3'd3,   
    WAIT_FOR_READ_SRAM_N_TH_DATA                = 3'd4,   
    WRITE_SRAM_ACCUMULATION            = 3'd5,   
    COMPUTE_COMPLETE              = 3'd6 } states;

states current_state, next_state;



always @(posedge clk) begin
// Synchronous active low reset.
if(!reset_n) begin
  // If reset stay in the idle state.
  dut_ready_reg <= 1'b1;
  current_state <= IDLE;
end else begin
  // if not in reset go to state 0 and read the 0th address.
  current_state <= next_state;
end
end


always @(*) begin : proc_next_state_fsm
  case (current_state)

    IDLE                    : begin
      if (dut_valid) begin
        set_dut_ready       = 1'b0;
        get_array_size      = 1'b0;
        read_addr_sel       = 2'b00;
        compute_accumulation= 1'b0;
        save_array_size     = 1'b0;
        write_enable_sel    = 1'b0;
        next_state          = READ_SRAM_ZERO_ADDR;
      end
      else begin
        set_dut_ready       = 1'b1;
        get_array_size      = 1'b0;
        read_addr_sel       = 2'b00;
        compute_accumulation= 1'b0;
        write_enable_sel    = 1'b0;
        save_array_size     = 1'b0;
        next_state          = IDLE;
      end
    end
  
    READ_SRAM_ZERO_ADDR  : begin
      set_dut_ready         = 1'b0;
      get_array_size        = 1'b1;
      read_addr_sel         = 2'b01;  // Increment the read addr
      compute_accumulation  = 1'b0;
      save_array_size       = 1'b0;
      write_enable_sel      = 1'b0;
      next_state            = READ_SRAM_FIRST_ARRAY_ELEMENT;
    end 

    READ_SRAM_FIRST_ARRAY_ELEMENT: begin
      set_dut_ready         = 1'b0;
      get_array_size        = 1'b0;
      read_addr_sel         = 2'b01;  // Increment the read addr
      compute_accumulation  = 1'b0;
      save_array_size       = 1'b1;
      write_enable_sel      = 1'b0;
      global_read_cycle_counter = matrixBRows * matrixBColumns;
      matrixBReadLimit      = matrixBColumns * matrixBRows;
      next_state            = READ_SRAM_2_N_ARRAY;    
    end

    READ_SRAM_2_N_ARRAY     : begin
      set_dut_ready         = 1'b0;
      get_array_size        = 1'b0;
      read_addr_sel         = 2'b01;  // Keep incrementing the read addr
      compute_accumulation  = 1'b1;
      save_array_size       = 1'b1;
      write_enable_sel      = 1'b0;
      next_state            = read_complete ? WAIT_FOR_READ_SRAM_N_TH_DATA : READ_SRAM_2_N_ARRAY;
    end 

    WAIT_FOR_READ_SRAM_N_TH_DATA : begin
      set_dut_ready         = 1'b0;
      get_array_size        = 1'b0;
      read_addr_sel         = 2'b10;  // Hold the address
      compute_accumulation  = 1'b1;
      save_array_size       = 1'b1;
      write_enable_sel      = 1'b0;
      next_state            = WRITE_SRAM_ACCUMULATION;    
    end

    WRITE_SRAM_ACCUMULATION : begin
      set_dut_ready         = 1'b0;
      get_array_size        = 1'b0;
      read_addr_sel         = 2'b10;  // Hold the address
      compute_accumulation  = 1'b0;
      save_array_size       = 1'b1;
      write_enable_sel      = 1'b1;
      next_state            = COMPUTE_COMPLETE;
    end

    COMPUTE_COMPLETE        : begin
      set_dut_ready         = 1'b1;
      get_array_size        = 1'b0;
      read_addr_sel         = 2'b00;  
      compute_accumulation  = 1'b0;
      save_array_size       = 1'b0;
      write_enable_sel      = 1'b0;
      next_state            = IDLE;      
    end

    default                 :  begin
      set_dut_ready         = 1'b1;
      get_array_size        = 1'b0;
      read_addr_sel         = 2'b00;  
      compute_accumulation  = 1'b0;
      save_array_size       = 1'b0;
      write_enable_sel      = 1'b0;      
      next_state            = IDLE;
    end
  endcase
end

always @(posedge clk) begin 
  if(!reset_n) begin
    compute_complete <= 0;
  end else begin
    compute_complete <= (dut_ready_reg) ? 1'b1 : 1'b0;
  end
end
  assign dut_ready = compute_complete;


always @(posedge clk) begin
  if(!reset_n) begin
    matrixAColumns  <= `SRAM_ADDR_WIDTH'b0;
    matrixARows     <= `SRAM_ADDR_WIDTH'b0;
    matrixBColumns  <= `SRAM_ADDR_WIDTH'b0;
    matrixBRows     <= `SRAM_ADDR_WIDTH'b0;
    matrix_A_read_counter    <= `SRAM_ADDR_WIDTH'b1;
    matrix_A_read_cycle_counter <= `SRAM_ADDR_WIDTH'b1;
    matrix_B_read_cycle_counter <= `SRAM_ADDR_WIDTH'b1;
    matrix_B_read_counter_1   <= `SRAM_ADDR_WIDTH'b1;
    matrix_B_read_counter_2   <= `SRAM_ADDR_WIDTH'b1;
    matrix_C_result_write_address_reg <= `SRAM_ADDR_WIDTH'b0;
    sram_result_write_address_reg <= `SRAM_ADDR_WIDTH'b0;
    matrix_A_address <= 1;
    matrix_A_row_counter <= 1;
    matrix_A_col_counter <= 1;
    matrix_B_row_repeat_counter <= 1;
  end else begin
    // If get_array_size is enabled in state, assign teh read data from sram to this register if not     
    matrixARows    <= get_array_size ? tb__dut__sram_input_read_data[31:16] : (save_array_size ? matrixARows : `SRAM_ADDR_WIDTH'b0);
    matrixAColumns <= get_array_size ? tb__dut__sram_input_read_data[15:0] : (save_array_size ? matrixAColumns : `SRAM_ADDR_WIDTH'b0);

    matrixBRows    <= get_array_size ? tb__dut__sram_weight_read_data[31:16] : (save_array_size ? matrixBRows : `SRAM_ADDR_WIDTH'b0);
    matrixBColumns <= get_array_size ? tb__dut__sram_weight_read_data[15:0] : (save_array_size ? matrixBColumns : `SRAM_ADDR_WIDTH'b0);
  end
end


// SRAM read address generator
always @(posedge clk) begin
    if (!reset_n) begin
      dut__tb__sram_input_read_address_reg  <= 0;
      dut__tb__sram_weight_read_address_reg  <= 0;
    end
    else begin

      case(read_addr_sel)

      2'b00 :begin 
                  dut__tb__sram_input_read_address_reg <= `SRAM_ADDR_WIDTH'b0;
                  dut__tb__sram_weight_read_address_reg <= `SRAM_ADDR_WIDTH'b0;
      end

      2'b01: begin
                  // Matrix A Address generator
        numOfReads <= numOfReads + 1;
        
      end

      2'b10: begin

        dut__tb__sram_input_read_address_reg <= dut__tb__sram_input_read_address_reg;
        dut__tb__sram_weight_read_address_reg <= dut__tb__sram_weight_read_address_reg;

      end


      default: begin
          dut__tb__sram_input_read_address_reg <= `SRAM_ADDR_WIDTH'b01;
          dut__tb__sram_weight_read_address_reg <= `SRAM_ADDR_WIDTH'b01;  
      end
      endcase

    end
        
end


always@(posedge clk) begin
if (!reset_n) begin
    dut__tb__sram_weight_read_address_reg <= `SRAM_DATA_WIDTH'b0;
    matrix_B_read_counter_1 <= `SRAM_DATA_WIDTH'b1;
    matrix_B_read_cycle_counter <= `SRAM_DATA_WIDTH'b1;
end
else if(read_addr_sel == 2'b01)begin
            // Matrix B Address generator
          if(matrix_B_read_cycle_counter <= matrixARows) begin
            if(matrix_B_read_counter_1 < matrixBReadLimit ) begin 
                    
              dut__tb__sram_weight_read_address_reg <= dut__tb__sram_weight_read_address_reg + `SRAM_DATA_WIDTH'b1;
              matrix_B_read_counter_1 <= matrix_B_read_counter_1 + `SRAM_DATA_WIDTH'b1;
              
            end else begin
              matrix_B_read_counter_1 <= `SRAM_DATA_WIDTH'b1;
              dut__tb__sram_weight_read_address_reg <= `SRAM_DATA_WIDTH'b1;
            end
          end else begin        
              matrix_B_read_cycle_counter <= matrix_B_read_cycle_counter + `SRAM_DATA_WIDTH'b1;   
          end
      end
end


assign dut__tb__sram_weight_read_address = dut__tb__sram_weight_read_address_reg;


always@(posedge clk) begin
if (!reset_n) begin
    dut__tb__sram_input_read_address_reg <= `SRAM_DATA_WIDTH'b0;
    matrix_A_col_counter <= `SRAM_DATA_WIDTH'b1;
    matrix_B_row_repeat_counter <= `SRAM_DATA_WIDTH'b1;
    sram_result_write_address_reg <= `SRAM_DATA_WIDTH'b0;
end
else if(read_addr_sel == 2'b01)begin
            // Repeat the same row Brow times
          if (matrix_B_row_repeat_counter <= matrixBRows) begin
        // Fetch the elements of the current row one at a time
            if (matrix_A_col_counter < matrixAColumns) begin
                // Assign the current read address to the SRAM input
                dut__tb__sram_input_read_address_reg <= (((matrix_A_row_counter - 1) * matrixAColumns) + matrix_A_col_counter);

                // Increment the column counter
                matrix_A_col_counter <= matrix_A_col_counter + 1;

                // Ensure write enable is low when fetching
                write_enable_sel <= 1'b0;

            end else begin
                // After fetching all columns in the row, reset column counter and increment repeat counter
                matrix_A_col_counter <= 1;  // Reset to 0 to start from the first column
                matrix_B_row_repeat_counter <= matrix_B_row_repeat_counter + 1;

                // Update SRAM input read address for the first column of the next fetch
                dut__tb__sram_input_read_address_reg <= (((matrix_A_row_counter - 1) * matrixAColumns) + matrix_A_col_counter);

                // Set write enable to high after fetching all columns
                write_enable_sel <= 1'b1;
                sram_result_write_address_reg <= sram_result_write_address_reg + 1;
            end
          end
      end
end

assign dut__tb__sram_input_read_address = dut__tb__sram_input_read_address_reg;



// READ N-elements in SRAM 
always @(posedge clk) begin : proc_read_completion
  if(!reset_n) begin
    
    read_complete <= 1'b0;
  end else begin
    read_complete <= (global_read_cycle_counter  == (matrixBReadLimit - 1)) ? 1'b1 : 1'b0;
  end
end

// SRAM write enable logic
always @(posedge clk) begin : proc_sram_write_enable_r
  if(!reset_n) begin
    dut__tb__sram_result_write_enable_reg <= 1'b0;
    dut__tb__sram_input_write_enable_reg <= 1'b0;
    dut__tb__sram_weight_write_enable_reg <= 1'b0;
  end else begin
    dut__tb__sram_result_write_enable_reg <= write_enable_sel ? 1'b1 : 1'b0;
  end
end

assign dut__tb__sram_result_write_enable = dut__tb__sram_result_write_enable_reg;
assign dut__tb__sram_input_write_enable = dut__tb__sram_input_write_enable_reg;
assign dut__tb__sram_weight_write_enable = dut__tb__sram_weight_write_enable_reg;


// SRAM write address logic
always @(posedge clk) begin : proc_sram_write_address_r
  if(!reset_n) begin
    dut__tb__sram_result_write_address_reg <= 1'b0;
  end else begin
    dut__tb__sram_result_write_address_reg <= (write_enable_sel) ? sram_result_write_address_reg : `SRAM_DATA_WIDTH'b0;  
  end
end

assign dut__tb__sram_result_write_address = dut__tb__sram_result_write_address_reg;
// SRAM write data logic
always @(posedge clk) begin : proc_sram_write_data_r
  if(!reset_n) begin
    dut__tb__sram_result_write_data_reg <= `SRAM_DATA_WIDTH'b0;
  end else begin
    dut__tb__sram_result_write_data_reg <= (write_enable_sel) ? sum_w : `SRAM_DATA_WIDTH'b0;
  end
end

assign dut__tb__sram_result_write_data = dut__tb__sram_result_write_data_reg;

// Accumulation logic 
always @(posedge clk) begin : proc_accumulation
  if(!reset_n) begin
    sum_r   <= `SRAM_DATA_WIDTH'b0;
  end else begin
    if (compute_accumulation) begin
      sum_r <= sum_w;
    end
    else begin
      sum_r <= `SRAM_DATA_WIDTH'b0;
    end
  end
end




// Floating-point multiply-accumulate instance
DW_fp_mac_inst FP_MAC (
  .inst_a(tb__dut__sram_input_read_data),
  .inst_b(tb__dut__sram_weight_read_data),
  .inst_c(sum_r),
  .inst_rnd(3'd0),
  .z_inst(sum_w),
  .status_inst()
);

endmodule


module DW_fp_mac_inst #(
  parameter inst_sig_width = 23,
  parameter inst_exp_width = 8,
  parameter inst_ieee_compliance = 0 // These need to be fixed to decrease error
) ( 
  input wire [inst_sig_width+inst_exp_width : 0] inst_a,
  input wire [inst_sig_width+inst_exp_width : 0] inst_b,
  input wire [inst_sig_width+inst_exp_width : 0] inst_c,
  input wire [2 : 0] inst_rnd,
  output wire [inst_sig_width+inst_exp_width : 0] z_inst,
  output wire [7 : 0] status_inst
);

  // Instance of DW_fp_mac
  DW_fp_mac #(inst_sig_width, inst_exp_width, inst_ieee_compliance) U1 (
    .a(inst_a),
    .b(inst_b),
    .c(inst_c),
    .rnd(inst_rnd),
    .z(z_inst),
    .status(status_inst) 
  );
endmodule